`define DBB_ADDR_START `NVDLA_MEM_ADDRESS_WIDTH'h8000_0000
`define DBB_MEM_SIZE (2**30-1)

//`define CVSRAM_ADDR_START `NVDLA_MEM_ADDRESS_WIDTH'h5000_0000
`define CVSRAM_ADDR_START `NVDLA_MEM_ADDRESS_WIDTH'h0000_0000
`define CVSRAM_MEM_SIZE (2**21-1)
